library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity galaga_cpu2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of galaga_cpu2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"00",X"91",X"C3",X"7C",X"05",X"FF",X"FF",X"87",X"30",X"05",X"24",X"C3",X"10",X"00",X"FF",
		X"85",X"6F",X"D0",X"24",X"C9",X"FF",X"FF",X"FF",X"77",X"23",X"10",X"FC",X"C9",X"23",X"06",X"16",
		X"23",X"00",X"19",X"F7",X"4B",X"00",X"23",X"F0",X"02",X"F0",X"5E",X"00",X"23",X"F0",X"24",X"FB",
		X"23",X"00",X"FF",X"FF",X"E9",X"FF",X"FF",X"FF",X"C3",X"13",X"05",X"BE",X"05",X"BF",X"05",X"D3",
		X"08",X"BE",X"05",X"F5",X"06",X"EE",X"05",X"BE",X"05",X"CA",X"0E",X"23",X"F0",X"26",X"23",X"14",
		X"13",X"FE",X"0D",X"0B",X"0A",X"08",X"06",X"04",X"03",X"01",X"23",X"FF",X"FF",X"FF",X"44",X"E4",
		X"18",X"FB",X"44",X"00",X"FF",X"FF",X"C9",X"23",X"08",X"08",X"23",X"03",X"1B",X"23",X"08",X"0F",
		X"23",X"16",X"15",X"F7",X"84",X"00",X"23",X"16",X"03",X"F0",X"97",X"00",X"23",X"16",X"19",X"FB",
		X"23",X"00",X"FF",X"FF",X"23",X"16",X"01",X"FE",X"0D",X"0C",X"0A",X"08",X"06",X"04",X"03",X"01",
		X"23",X"FC",X"30",X"23",X"00",X"FF",X"FF",X"44",X"27",X"0E",X"FB",X"44",X"00",X"FF",X"FF",X"33",
		X"06",X"18",X"23",X"00",X"18",X"F7",X"B6",X"00",X"23",X"F0",X"08",X"F0",X"CC",X"00",X"23",X"F0",
		X"20",X"FB",X"23",X"00",X"FF",X"FF",X"23",X"F0",X"20",X"23",X"10",X"0D",X"FE",X"1A",X"18",X"15",
		X"10",X"0C",X"08",X"05",X"03",X"23",X"FE",X"30",X"23",X"00",X"FF",X"FF",X"33",X"E0",X"10",X"FB",
		X"44",X"00",X"FF",X"FF",X"23",X"03",X"18",X"33",X"04",X"10",X"23",X"08",X"0A",X"44",X"16",X"12",
		X"F7",X"60",X"01",X"44",X"16",X"03",X"F0",X"73",X"01",X"44",X"16",X"1D",X"FB",X"23",X"00",X"FF",
		X"FF",X"12",X"18",X"17",X"12",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"14",X"06",X"14",X"0C",X"14",X"08",X"14",X"0A",X"1C",X"00",X"1C",X"12",X"1E",X"00",X"1E",X"12",
		X"1C",X"02",X"1C",X"10",X"1E",X"02",X"1E",X"10",X"1C",X"04",X"1C",X"0E",X"1E",X"04",X"1E",X"0E",
		X"1C",X"06",X"1C",X"0C",X"1E",X"06",X"1E",X"0C",X"1C",X"08",X"1C",X"0A",X"1E",X"08",X"1E",X"0A",
		X"16",X"06",X"16",X"0C",X"16",X"08",X"16",X"0A",X"18",X"00",X"18",X"12",X"1A",X"00",X"1A",X"12",
		X"18",X"02",X"18",X"10",X"1A",X"02",X"1A",X"10",X"18",X"04",X"18",X"0E",X"1A",X"04",X"1A",X"0E",
		X"18",X"06",X"18",X"0C",X"1A",X"06",X"1A",X"0C",X"18",X"08",X"18",X"0A",X"1A",X"08",X"1A",X"0A",
		X"44",X"16",X"06",X"FE",X"0C",X"0B",X"0A",X"08",X"06",X"04",X"02",X"01",X"23",X"FE",X"30",X"23",
		X"00",X"FF",X"FF",X"66",X"20",X"14",X"FB",X"44",X"00",X"FF",X"FF",X"23",X"06",X"18",X"23",X"00",
		X"18",X"F7",X"92",X"01",X"44",X"F0",X"08",X"F0",X"A8",X"01",X"44",X"F0",X"20",X"FB",X"23",X"00",
		X"FF",X"FF",X"44",X"F0",X"26",X"23",X"10",X"0B",X"FE",X"22",X"20",X"1E",X"1B",X"18",X"15",X"12",
		X"10",X"23",X"FE",X"30",X"23",X"00",X"FF",X"FF",X"66",X"E0",X"10",X"FB",X"44",X"00",X"FF",X"FF",
		X"23",X"03",X"20",X"23",X"08",X"0F",X"23",X"16",X"12",X"F7",X"CA",X"01",X"23",X"16",X"03",X"F0",
		X"E0",X"01",X"23",X"16",X"1D",X"FB",X"23",X"00",X"FF",X"FF",X"23",X"16",X"01",X"FE",X"0D",X"0C",
		X"0B",X"09",X"07",X"05",X"03",X"02",X"23",X"02",X"20",X"23",X"FC",X"12",X"23",X"00",X"FF",X"FF",
		X"44",X"20",X"14",X"FB",X"44",X"00",X"FF",X"FF",X"23",X"00",X"10",X"23",X"01",X"40",X"22",X"0C",
		X"37",X"23",X"00",X"FF",X"FF",X"23",X"02",X"3A",X"23",X"10",X"09",X"23",X"00",X"18",X"23",X"20",
		X"10",X"23",X"00",X"18",X"23",X"20",X"0D",X"23",X"00",X"FF",X"FF",X"23",X"00",X"10",X"23",X"01",
		X"30",X"00",X"40",X"08",X"23",X"FF",X"30",X"23",X"00",X"FF",X"FF",X"23",X"00",X"30",X"23",X"05",
		X"80",X"23",X"05",X"4C",X"23",X"04",X"01",X"23",X"00",X"50",X"FF",X"23",X"00",X"28",X"23",X"06",
		X"1D",X"23",X"00",X"11",X"00",X"40",X"08",X"23",X"00",X"11",X"23",X"FA",X"1D",X"23",X"00",X"50",
		X"FF",X"23",X"00",X"21",X"00",X"20",X"10",X"23",X"F8",X"20",X"23",X"FF",X"20",X"23",X"F8",X"1B",
		X"23",X"E8",X"0B",X"23",X"00",X"21",X"00",X"20",X"08",X"23",X"00",X"42",X"FF",X"23",X"00",X"08",
		X"00",X"20",X"08",X"23",X"F0",X"20",X"23",X"10",X"20",X"23",X"F0",X"40",X"23",X"10",X"20",X"23",
		X"F0",X"20",X"00",X"20",X"08",X"23",X"00",X"30",X"FF",X"23",X"10",X"0C",X"23",X"00",X"20",X"23",
		X"E8",X"10",X"23",X"F4",X"10",X"23",X"E8",X"10",X"23",X"F4",X"32",X"23",X"E8",X"10",X"23",X"F4",
		X"32",X"23",X"E8",X"10",X"23",X"F4",X"10",X"23",X"E8",X"0E",X"23",X"02",X"30",X"FF",X"23",X"F1",
		X"08",X"23",X"00",X"10",X"23",X"05",X"3C",X"23",X"07",X"42",X"23",X"0A",X"40",X"23",X"10",X"2D",
		X"23",X"20",X"19",X"00",X"FC",X"14",X"23",X"02",X"4A",X"FF",X"23",X"04",X"20",X"23",X"00",X"16",
		X"23",X"F0",X"30",X"23",X"00",X"12",X"23",X"10",X"30",X"23",X"00",X"12",X"23",X"10",X"30",X"23",
		X"00",X"16",X"23",X"04",X"20",X"23",X"00",X"10",X"FF",X"23",X"00",X"15",X"00",X"20",X"08",X"23",
		X"00",X"11",X"00",X"E0",X"08",X"23",X"00",X"18",X"00",X"20",X"08",X"23",X"00",X"13",X"00",X"E0",
		X"08",X"23",X"00",X"1F",X"00",X"20",X"08",X"23",X"00",X"30",X"FF",X"23",X"02",X"0E",X"23",X"00",
		X"34",X"23",X"12",X"19",X"23",X"00",X"20",X"23",X"E0",X"0E",X"23",X"00",X"12",X"23",X"20",X"0E",
		X"23",X"00",X"0C",X"23",X"E0",X"0E",X"23",X"1B",X"08",X"23",X"00",X"10",X"FF",X"23",X"00",X"0D",
		X"00",X"C0",X"04",X"23",X"00",X"21",X"00",X"40",X"06",X"23",X"00",X"51",X"00",X"C0",X"06",X"23",
		X"00",X"73",X"FF",X"23",X"08",X"20",X"23",X"00",X"16",X"23",X"E0",X"0C",X"23",X"02",X"0B",X"23",
		X"11",X"0C",X"23",X"02",X"0B",X"23",X"E0",X"0C",X"23",X"00",X"16",X"23",X"08",X"20",X"FF",X"12",
		X"18",X"1E",X"12",X"00",X"34",X"12",X"FB",X"26",X"12",X"00",X"02",X"FC",X"2E",X"12",X"FA",X"3C",
		X"FA",X"9E",X"03",X"12",X"F8",X"10",X"12",X"FA",X"5C",X"12",X"00",X"23",X"F8",X"F9",X"EF",X"7C",
		X"03",X"F6",X"AB",X"12",X"01",X"28",X"12",X"0A",X"18",X"FD",X"52",X"03",X"F6",X"B0",X"23",X"08",
		X"1E",X"23",X"00",X"19",X"23",X"F8",X"16",X"23",X"00",X"02",X"FC",X"30",X"23",X"F7",X"26",X"FA",
		X"9E",X"03",X"23",X"F0",X"0A",X"23",X"F5",X"31",X"23",X"00",X"10",X"FD",X"6C",X"03",X"12",X"F8",
		X"10",X"12",X"00",X"40",X"FB",X"12",X"00",X"FF",X"FF",X"12",X"18",X"1D",X"12",X"00",X"28",X"12",
		X"FA",X"02",X"F3",X"3F",X"3B",X"36",X"32",X"28",X"26",X"24",X"22",X"12",X"04",X"30",X"12",X"FC",
		X"30",X"12",X"00",X"18",X"F8",X"F9",X"FA",X"0C",X"04",X"EF",X"D7",X"03",X"F6",X"B0",X"12",X"01",
		X"28",X"12",X"0A",X"15",X"FD",X"AC",X"03",X"F6",X"C0",X"23",X"08",X"10",X"23",X"00",X"23",X"23",
		X"F8",X"0F",X"23",X"00",X"48",X"F8",X"F9",X"FA",X"0C",X"04",X"F6",X"B0",X"23",X"08",X"20",X"23",
		X"00",X"08",X"23",X"F8",X"02",X"F3",X"34",X"31",X"2D",X"29",X"22",X"26",X"1F",X"18",X"23",X"08",
		X"18",X"23",X"F8",X"18",X"23",X"00",X"10",X"F8",X"F9",X"FD",X"CC",X"03",X"FB",X"12",X"00",X"FF",
		X"FF",X"12",X"18",X"14",X"12",X"03",X"2A",X"12",X"10",X"40",X"12",X"01",X"20",X"12",X"FE",X"71",
		X"F9",X"F1",X"FA",X"0C",X"04",X"EF",X"30",X"04",X"F6",X"AB",X"12",X"02",X"20",X"FD",X"14",X"04",
		X"F6",X"B0",X"23",X"04",X"1A",X"23",X"03",X"1D",X"23",X"1A",X"25",X"23",X"03",X"10",X"23",X"FD",
		X"48",X"FD",X"20",X"04",X"12",X"18",X"14",X"12",X"03",X"2A",X"12",X"10",X"40",X"12",X"01",X"20",
		X"12",X"FE",X"78",X"FF",X"12",X"18",X"14",X"F4",X"12",X"00",X"04",X"FC",X"48",X"00",X"FC",X"FF",
		X"23",X"00",X"30",X"F8",X"F9",X"FA",X"0C",X"04",X"FD",X"25",X"04",X"12",X"18",X"14",X"FB",X"12",
		X"00",X"FF",X"FF",X"12",X"18",X"1E",X"12",X"00",X"08",X"F2",X"99",X"04",X"00",X"00",X"0A",X"F2",
		X"99",X"04",X"00",X"00",X"0A",X"12",X"00",X"2C",X"12",X"FB",X"26",X"12",X"00",X"02",X"FC",X"2E",
		X"12",X"FA",X"3C",X"FA",X"9E",X"03",X"FD",X"63",X"03",X"12",X"00",X"2C",X"12",X"FB",X"26",X"12",
		X"00",X"02",X"FC",X"2E",X"12",X"FA",X"18",X"12",X"00",X"10",X"FF",X"12",X"18",X"13",X"F2",X"C6",
		X"04",X"00",X"00",X"08",X"F2",X"CF",X"04",X"00",X"00",X"08",X"12",X"18",X"0B",X"12",X"00",X"34",
		X"12",X"FB",X"26",X"FD",X"58",X"03",X"12",X"00",X"10",X"12",X"18",X"0B",X"FD",X"D8",X"04",X"12",
		X"00",X"08",X"12",X"18",X"0B",X"12",X"00",X"06",X"12",X"00",X"22",X"12",X"FB",X"26",X"12",X"00",
		X"02",X"FC",X"2E",X"12",X"FA",X"18",X"12",X"00",X"20",X"FF",X"12",X"18",X"1E",X"12",X"00",X"14",
		X"F2",X"02",X"05",X"12",X"00",X"08",X"F2",X"02",X"05",X"12",X"00",X"18",X"12",X"FB",X"26",X"FD",
		X"58",X"03",X"12",X"E2",X"01",X"F3",X"08",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"F5",X"23",
		X"00",X"48",X"FF",X"AF",X"32",X"21",X"68",X"3A",X"04",X"68",X"E6",X"02",X"CA",X"75",X"05",X"3A",
		X"A0",X"92",X"3C",X"32",X"A0",X"92",X"2A",X"A1",X"92",X"E6",X"1F",X"3D",X"28",X"08",X"3C",X"20",
		X"06",X"7C",X"F6",X"01",X"67",X"2C",X"24",X"22",X"A1",X"92",X"3A",X"C7",X"99",X"5F",X"3A",X"A7",
		X"92",X"BB",X"CB",X"10",X"3A",X"15",X"90",X"A0",X"E6",X"01",X"32",X"AA",X"92",X"0E",X"00",X"21",
		X"20",X"90",X"79",X"85",X"6F",X"7E",X"A7",X"20",X"03",X"0C",X"18",X"F3",X"47",X"21",X"3B",X"00",
		X"79",X"CB",X"27",X"85",X"6F",X"5E",X"23",X"56",X"EB",X"C5",X"CD",X"34",X"00",X"C1",X"78",X"81",
		X"4F",X"E6",X"F8",X"28",X"DA",X"3E",X"01",X"32",X"21",X"68",X"FB",X"C9",X"11",X"00",X"91",X"1A",
		X"A7",X"20",X"FC",X"67",X"6F",X"01",X"10",X"00",X"86",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"FE",
		X"FF",X"28",X"02",X"3E",X"11",X"12",X"1A",X"A7",X"20",X"FC",X"ED",X"56",X"AF",X"32",X"E0",X"89",
		X"21",X"B7",X"05",X"11",X"21",X"90",X"01",X"07",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"21",X"68",
		X"FB",X"31",X"00",X"91",X"C3",X"B1",X"05",X"01",X"01",X"00",X"01",X"01",X"00",X"0A",X"C9",X"3E",
		X"01",X"32",X"D7",X"92",X"21",X"00",X"8B",X"11",X"80",X"8B",X"01",X"40",X"00",X"ED",X"B0",X"21",
		X"00",X"93",X"11",X"80",X"93",X"0E",X"40",X"ED",X"B0",X"21",X"00",X"9B",X"11",X"80",X"9B",X"0E",
		X"40",X"ED",X"B0",X"AF",X"32",X"D7",X"92",X"3A",X"D6",X"92",X"3D",X"28",X"FA",X"C9",X"3A",X"14",
		X"90",X"A7",X"C8",X"32",X"17",X"92",X"3A",X"27",X"98",X"A7",X"28",X"17",X"21",X"60",X"93",X"7E",
		X"A7",X"28",X"10",X"CD",X"81",X"06",X"3A",X"BF",X"99",X"A7",X"28",X"07",X"CD",X"49",X"06",X"AF",
		X"32",X"2B",X"98",X"21",X"62",X"93",X"7E",X"A7",X"C8",X"CD",X"81",X"06",X"3A",X"BF",X"99",X"A7",
		X"C8",X"3A",X"27",X"98",X"A7",X"28",X"12",X"AF",X"32",X"2B",X"98",X"3A",X"60",X"93",X"32",X"62",
		X"93",X"3A",X"E2",X"93",X"21",X"E0",X"93",X"18",X"16",X"AF",X"32",X"14",X"90",X"32",X"15",X"90",
		X"32",X"25",X"90",X"32",X"B9",X"99",X"32",X"17",X"92",X"EB",X"26",X"93",X"CB",X"FD",X"7E",X"D6",
		X"08",X"CB",X"BD",X"77",X"2C",X"7E",X"D6",X"08",X"77",X"26",X"8B",X"36",X"0B",X"2D",X"36",X"20",
		X"26",X"88",X"36",X"08",X"2C",X"36",X"0F",X"2D",X"26",X"9B",X"36",X"0C",X"AF",X"32",X"27",X"98",
		X"3A",X"01",X"92",X"3D",X"32",X"B9",X"9A",X"3A",X"17",X"92",X"A7",X"C0",X"3C",X"32",X"13",X"92",
		X"C9",X"AF",X"32",X"BF",X"99",X"26",X"88",X"7E",X"26",X"93",X"FE",X"08",X"C8",X"7E",X"DD",X"6F",
		X"2C",X"46",X"26",X"9B",X"7E",X"0F",X"CB",X"18",X"DD",X"60",X"2D",X"5D",X"3A",X"08",X"90",X"A7",
		X"28",X"06",X"2E",X"38",X"06",X"04",X"18",X"04",X"2E",X"00",X"06",X"30",X"CD",X"B7",X"06",X"2E",
		X"68",X"06",X"08",X"CD",X"B7",X"06",X"C9",X"26",X"92",X"7E",X"26",X"88",X"B6",X"07",X"38",X"30",
		X"7E",X"E6",X"FE",X"FE",X"04",X"28",X"29",X"26",X"93",X"7E",X"A7",X"28",X"23",X"DD",X"95",X"D6",
		X"07",X"C6",X"0D",X"30",X"1B",X"2C",X"7E",X"26",X"9B",X"4E",X"2D",X"CB",X"09",X"1F",X"DD",X"94",
		X"D6",X"04",X"C6",X"07",X"30",X"0A",X"3E",X"01",X"32",X"BF",X"99",X"B7",X"08",X"C3",X"C2",X"07",
		X"2C",X"2C",X"10",X"C3",X"C9",X"11",X"A4",X"92",X"21",X"64",X"93",X"CD",X"04",X"07",X"11",X"A5",
		X"92",X"21",X"66",X"93",X"7E",X"A7",X"C8",X"1A",X"47",X"E6",X"07",X"08",X"3E",X"06",X"CB",X"78",
		X"28",X"01",X"08",X"CB",X"70",X"28",X"02",X"ED",X"44",X"86",X"77",X"FE",X"F0",X"30",X"44",X"DD",
		X"6F",X"2C",X"08",X"CB",X"68",X"28",X"02",X"ED",X"44",X"4F",X"86",X"77",X"1F",X"A9",X"26",X"9B",
		X"07",X"30",X"05",X"CB",X"0E",X"3F",X"CB",X"16",X"4E",X"26",X"93",X"7E",X"CB",X"09",X"1F",X"DD",
		X"67",X"FE",X"14",X"38",X"1B",X"FE",X"9C",X"30",X"17",X"5D",X"3A",X"1D",X"90",X"A7",X"28",X"07",
		X"21",X"08",X"93",X"06",X"2C",X"18",X"05",X"21",X"00",X"93",X"06",X"30",X"CD",X"6A",X"07",X"C9",
		X"2D",X"26",X"93",X"36",X"00",X"26",X"9B",X"36",X"00",X"C9",X"26",X"92",X"7E",X"26",X"88",X"B6",
		X"07",X"38",X"41",X"7E",X"4F",X"E6",X"FE",X"FE",X"04",X"28",X"39",X"2C",X"26",X"9B",X"56",X"26",
		X"93",X"7E",X"CB",X"0A",X"1F",X"2D",X"DD",X"94",X"D6",X"03",X"C6",X"06",X"30",X"26",X"79",X"3D",
		X"E6",X"FE",X"08",X"3A",X"27",X"98",X"A7",X"7E",X"20",X"0A",X"DD",X"95",X"D6",X"06",X"C6",X"0B",
		X"38",X"17",X"18",X"10",X"DD",X"95",X"D6",X"14",X"C6",X"0B",X"38",X"0D",X"C6",X"04",X"38",X"04",
		X"C6",X"0B",X"38",X"05",X"2C",X"2C",X"10",X"B2",X"C9",X"7D",X"2A",X"44",X"98",X"23",X"22",X"44",
		X"98",X"6F",X"16",X"93",X"AF",X"12",X"16",X"9B",X"12",X"2C",X"26",X"8B",X"7E",X"4F",X"A7",X"CA",
		X"CA",X"08",X"2D",X"FE",X"0B",X"28",X"3E",X"08",X"20",X"44",X"08",X"26",X"92",X"36",X"81",X"3A",
		X"28",X"98",X"95",X"20",X"07",X"32",X"2B",X"98",X"3C",X"32",X"28",X"98",X"E5",X"79",X"FE",X"07",
		X"20",X"03",X"3D",X"18",X"03",X"3D",X"E6",X"03",X"21",X"A1",X"9A",X"D7",X"36",X"01",X"79",X"FE",
		X"07",X"20",X"05",X"21",X"2B",X"98",X"36",X"00",X"21",X"90",X"92",X"D7",X"34",X"08",X"28",X"01",
		X"34",X"E1",X"C3",X"B4",X"07",X"26",X"93",X"36",X"00",X"26",X"88",X"36",X"80",X"C9",X"26",X"88",
		X"E5",X"08",X"2C",X"7E",X"26",X"91",X"C6",X"13",X"6F",X"36",X"00",X"21",X"88",X"92",X"34",X"21",
		X"A8",X"92",X"35",X"E1",X"20",X"13",X"26",X"92",X"3A",X"85",X"92",X"77",X"3A",X"84",X"92",X"67",
		X"3A",X"9F",X"92",X"84",X"32",X"9F",X"92",X"18",X"96",X"79",X"FE",X"07",X"20",X"04",X"16",X"B8",
		X"18",X"5E",X"3A",X"2D",X"98",X"BD",X"CA",X"B6",X"08",X"7D",X"E6",X"38",X"FE",X"38",X"CA",X"B6",
		X"08",X"79",X"FE",X"01",X"C2",X"DB",X"07",X"D5",X"7D",X"E6",X"07",X"5F",X"16",X"88",X"1A",X"FE",
		X"09",X"20",X"26",X"E5",X"EB",X"2C",X"7E",X"C6",X"13",X"5F",X"16",X"91",X"AF",X"12",X"26",X"8B",
		X"36",X"09",X"2D",X"7D",X"32",X"28",X"98",X"26",X"88",X"AF",X"77",X"32",X"8B",X"92",X"3C",X"32",
		X"1D",X"90",X"32",X"8D",X"92",X"32",X"B1",X"9A",X"E1",X"D1",X"E5",X"3E",X"06",X"32",X"AD",X"92",
		X"7D",X"E6",X"07",X"21",X"30",X"98",X"D7",X"7E",X"2C",X"56",X"21",X"9F",X"92",X"86",X"77",X"E1",
		X"26",X"92",X"72",X"C3",X"DF",X"07",X"E5",X"21",X"B0",X"99",X"35",X"E1",X"C2",X"DB",X"07",X"3A",
		X"B2",X"99",X"57",X"3A",X"B1",X"99",X"E5",X"C3",X"AA",X"08",X"3C",X"77",X"32",X"A4",X"9A",X"2D",
		X"C3",X"B4",X"07",X"DD",X"21",X"00",X"91",X"3E",X"0C",X"32",X"89",X"92",X"21",X"86",X"92",X"7E",
		X"36",X"00",X"23",X"77",X"DD",X"CB",X"13",X"46",X"CA",X"FA",X"0D",X"21",X"86",X"92",X"34",X"DD",
		X"6E",X"10",X"26",X"88",X"7E",X"FE",X"03",X"28",X"09",X"FE",X"09",X"28",X"05",X"FE",X"07",X"C2",
		X"48",X"0E",X"DD",X"35",X"0D",X"C2",X"00",X"0C",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"7E",X"FE",
		X"EF",X"DA",X"D7",X"0B",X"E5",X"2F",X"21",X"20",X"09",X"CF",X"7E",X"23",X"66",X"6F",X"E3",X"C9",
		X"48",X"0E",X"11",X"0B",X"41",X"0B",X"49",X"0B",X"9B",X"0A",X"CC",X"0B",X"5A",X"0B",X"82",X"0B",
		X"93",X"0B",X"A3",X"0B",X"42",X"09",X"50",X"0A",X"FE",X"09",X"7B",X"09",X"68",X"09",X"55",X"09",
		X"4E",X"09",X"DD",X"5E",X"10",X"16",X"88",X"3E",X"03",X"12",X"23",X"C3",X"0E",X"09",X"3A",X"C9",
		X"99",X"A7",X"C3",X"59",X"09",X"3A",X"C8",X"99",X"A7",X"28",X"08",X"23",X"7E",X"23",X"66",X"6F",
		X"C3",X"87",X"0B",X"23",X"23",X"C3",X"86",X"0B",X"DD",X"5E",X"10",X"16",X"01",X"1A",X"5F",X"16",
		X"99",X"1C",X"1A",X"C6",X"20",X"DD",X"77",X"01",X"C3",X"86",X"0B",X"E5",X"DD",X"5E",X"10",X"21",
		X"38",X"88",X"06",X"04",X"7E",X"07",X"38",X"07",X"2C",X"2C",X"10",X"F8",X"C3",X"FA",X"09",X"26",
		X"8B",X"54",X"1A",X"77",X"2C",X"1C",X"1A",X"77",X"2D",X"7D",X"08",X"21",X"EF",X"91",X"11",X"EC",
		X"FF",X"06",X"0C",X"7E",X"E6",X"01",X"28",X"06",X"19",X"10",X"F8",X"C3",X"FA",X"09",X"19",X"23",
		X"DD",X"7E",X"00",X"DD",X"5D",X"DD",X"54",X"EB",X"FD",X"6B",X"FD",X"62",X"01",X"06",X"00",X"ED",
		X"B0",X"0E",X"06",X"09",X"EB",X"19",X"EB",X"0E",X"04",X"ED",X"B0",X"DD",X"7E",X"13",X"FD",X"77",
		X"13",X"E1",X"23",X"7E",X"FD",X"77",X"08",X"23",X"7E",X"FD",X"77",X"09",X"FD",X"36",X"0A",X"01",
		X"FD",X"36",X"0B",X"02",X"FD",X"36",X"0D",X"01",X"08",X"FD",X"77",X"10",X"5F",X"16",X"88",X"3E",
		X"09",X"12",X"1C",X"FD",X"7D",X"12",X"23",X"C3",X"0E",X"09",X"E1",X"C3",X"9D",X"0B",X"E5",X"EB",
		X"3A",X"15",X"92",X"4F",X"3A",X"62",X"93",X"FE",X"1E",X"30",X"02",X"3E",X"1E",X"FE",X"D1",X"38",
		X"02",X"3E",X"D1",X"CB",X"41",X"28",X"04",X"C6",X"0E",X"ED",X"44",X"CB",X"3F",X"DD",X"96",X"03",
		X"1F",X"DD",X"CB",X"13",X"7E",X"28",X"02",X"ED",X"44",X"C6",X"18",X"F2",X"2F",X"0A",X"AF",X"FE",
		X"30",X"38",X"02",X"3E",X"2F",X"67",X"3E",X"06",X"CD",X"A9",X"0E",X"7C",X"3C",X"EB",X"D7",X"7E",
		X"DD",X"77",X"0D",X"E1",X"3E",X"09",X"D7",X"DD",X"75",X"08",X"DD",X"74",X"09",X"C3",X"FA",X"0B",
		X"E5",X"3A",X"15",X"92",X"4F",X"3A",X"62",X"93",X"C6",X"03",X"E6",X"F8",X"3C",X"FE",X"29",X"30",
		X"02",X"3E",X"29",X"FE",X"CA",X"38",X"02",X"3E",X"C9",X"CB",X"41",X"28",X"03",X"C6",X"0D",X"2F",
		X"32",X"8A",X"92",X"CB",X"3F",X"5F",X"16",X"48",X"DD",X"66",X"01",X"DD",X"6E",X"03",X"CD",X"5A",
		X"0E",X"CB",X"3C",X"CB",X"1D",X"DD",X"75",X"04",X"DD",X"74",X"05",X"AF",X"32",X"8B",X"92",X"3C",
		X"32",X"19",X"90",X"DD",X"7D",X"32",X"29",X"98",X"C3",X"0C",X"0B",X"E5",X"DD",X"6E",X"10",X"26",
		X"88",X"36",X"09",X"26",X"01",X"4E",X"2C",X"6E",X"26",X"99",X"46",X"2C",X"5E",X"69",X"4E",X"2C",
		X"56",X"CB",X"3B",X"D5",X"DD",X"70",X"11",X"DD",X"71",X"12",X"3A",X"15",X"92",X"A7",X"28",X"08",
		X"78",X"ED",X"44",X"47",X"79",X"ED",X"44",X"4F",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"51",X"1E",
		X"00",X"CB",X"2A",X"CB",X"1B",X"19",X"DD",X"75",X"00",X"DD",X"74",X"01",X"5C",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"0E",X"00",X"CB",X"28",X"CB",X"19",X"ED",X"42",X"DD",X"75",X"02",X"DD",X"74",
		X"03",X"6C",X"63",X"4A",X"D1",X"CD",X"5A",X"0E",X"CB",X"3C",X"CB",X"1D",X"DD",X"75",X"04",X"DD",
		X"74",X"05",X"DD",X"72",X"06",X"DD",X"73",X"07",X"DD",X"CB",X"13",X"F6",X"E1",X"23",X"C3",X"0E",
		X"09",X"E5",X"EB",X"3A",X"15",X"92",X"0F",X"DD",X"46",X"13",X"A8",X"07",X"3A",X"E2",X"93",X"3C",
		X"3D",X"20",X"02",X"3E",X"80",X"38",X"04",X"ED",X"44",X"C6",X"F2",X"C6",X"0E",X"67",X"3E",X"1E",
		X"CD",X"A9",X"0E",X"7C",X"EB",X"D7",X"7E",X"DD",X"77",X"0D",X"E1",X"3E",X"09",X"D7",X"C3",X"FA",
		X"0B",X"23",X"5E",X"23",X"56",X"EB",X"C3",X"0E",X"09",X"23",X"5E",X"23",X"DD",X"73",X"06",X"DD",
		X"36",X"07",X"00",X"DD",X"CB",X"13",X"EE",X"C3",X"FA",X"0B",X"3A",X"15",X"92",X"4F",X"DD",X"5E",
		X"10",X"1C",X"16",X"01",X"1A",X"5F",X"16",X"98",X"1A",X"CB",X"41",X"28",X"04",X"C6",X"0E",X"ED",
		X"44",X"CB",X"3F",X"DD",X"77",X"03",X"3A",X"AA",X"92",X"A7",X"CA",X"86",X"0B",X"32",X"B3",X"9A",
		X"18",X"04",X"DD",X"36",X"01",X"9C",X"23",X"DD",X"75",X"08",X"DD",X"74",X"09",X"DD",X"34",X"0D",
		X"C3",X"FA",X"0D",X"DD",X"7E",X"10",X"E6",X"38",X"FE",X"38",X"CA",X"41",X"0B",X"23",X"23",X"23",
		X"C3",X"0E",X"09",X"23",X"7E",X"DD",X"CB",X"13",X"7E",X"28",X"04",X"C6",X"80",X"ED",X"44",X"0E",
		X"00",X"CB",X"27",X"CB",X"11",X"CB",X"27",X"CB",X"11",X"DD",X"77",X"04",X"DD",X"71",X"05",X"DD",
		X"36",X"0E",X"1E",X"3A",X"C8",X"92",X"DD",X"77",X"0F",X"C3",X"86",X"0B",X"3A",X"AA",X"92",X"4F",
		X"3A",X"1D",X"90",X"3D",X"A1",X"18",X"C3",X"4F",X"E6",X"0F",X"DD",X"77",X"0A",X"79",X"07",X"07",
		X"07",X"07",X"E6",X"0F",X"23",X"DD",X"77",X"0B",X"7E",X"23",X"DD",X"CB",X"13",X"7E",X"28",X"02",
		X"ED",X"44",X"DD",X"77",X"0C",X"7E",X"23",X"DD",X"77",X"0D",X"DD",X"75",X"08",X"DD",X"74",X"09",
		X"DD",X"CB",X"13",X"76",X"28",X"22",X"DD",X"7E",X"01",X"DD",X"96",X"06",X"28",X"08",X"F2",X"13",
		X"0C",X"ED",X"44",X"3D",X"20",X"12",X"DD",X"7E",X"03",X"DD",X"96",X"07",X"CA",X"07",X"0E",X"F2",
		X"24",X"0C",X"ED",X"44",X"3D",X"CA",X"07",X"0E",X"DD",X"CB",X"13",X"6E",X"28",X"13",X"DD",X"7E",
		X"01",X"DD",X"96",X"06",X"28",X"03",X"3C",X"20",X"08",X"DD",X"36",X"0D",X"01",X"DD",X"CB",X"13",
		X"AE",X"DD",X"46",X"0C",X"DD",X"7E",X"04",X"5F",X"80",X"DD",X"77",X"04",X"DD",X"56",X"05",X"2E",
		X"01",X"CB",X"78",X"28",X"02",X"2E",X"FF",X"1F",X"A8",X"7A",X"F2",X"5E",X"0C",X"85",X"DD",X"77",
		X"05",X"7B",X"4A",X"CB",X"41",X"28",X"01",X"2F",X"C6",X"15",X"30",X"04",X"06",X"06",X"18",X"0C",
		X"CB",X"3F",X"47",X"CB",X"38",X"80",X"07",X"07",X"07",X"E6",X"07",X"47",X"26",X"8B",X"DD",X"6E",
		X"10",X"7E",X"E6",X"F8",X"B0",X"77",X"26",X"9B",X"79",X"CB",X"09",X"A9",X"3C",X"CB",X"09",X"17",
		X"E6",X"03",X"77",X"3A",X"A0",X"92",X"E6",X"01",X"28",X"05",X"DD",X"7E",X"0A",X"18",X"03",X"DD",
		X"7E",X"0B",X"A7",X"CA",X"FE",X"0C",X"E5",X"DD",X"E5",X"E1",X"47",X"7A",X"E6",X"03",X"57",X"CB",
		X"03",X"CB",X"12",X"D5",X"AA",X"0F",X"38",X"02",X"2C",X"2C",X"14",X"CB",X"52",X"78",X"28",X"02",
		X"ED",X"44",X"4F",X"CB",X"29",X"30",X"04",X"7E",X"C6",X"80",X"77",X"2C",X"7E",X"89",X"77",X"2D",
		X"EB",X"7B",X"EE",X"02",X"5F",X"E1",X"CB",X"3D",X"30",X"04",X"7D",X"EE",X"7F",X"6F",X"78",X"44",
		X"26",X"00",X"CD",X"96",X"0E",X"78",X"EE",X"02",X"3D",X"CB",X"57",X"28",X"08",X"44",X"4D",X"21",
		X"00",X"00",X"A7",X"ED",X"42",X"EB",X"7B",X"86",X"77",X"2C",X"7A",X"8E",X"77",X"E1",X"3A",X"15",
		X"92",X"4F",X"26",X"93",X"DD",X"56",X"03",X"3E",X"7F",X"DD",X"BE",X"02",X"7A",X"17",X"CB",X"41",
		X"28",X"03",X"C6",X"0D",X"2F",X"DD",X"CB",X"13",X"76",X"28",X"03",X"DD",X"86",X"11",X"77",X"2C",
		X"DD",X"46",X"01",X"3E",X"7F",X"DD",X"BE",X"00",X"CB",X"13",X"78",X"CB",X"41",X"20",X"04",X"C6",
		X"4F",X"2F",X"1D",X"CB",X"1B",X"17",X"CB",X"13",X"DD",X"CB",X"13",X"76",X"28",X"0D",X"DD",X"86",
		X"12",X"57",X"1F",X"DD",X"AE",X"12",X"07",X"7A",X"30",X"01",X"1C",X"77",X"26",X"9B",X"CB",X"0E",
		X"CB",X"0B",X"CB",X"16",X"DD",X"35",X"0E",X"C2",X"FA",X"0D",X"DD",X"CB",X"0F",X"3E",X"D2",X"F4",
		X"0D",X"DD",X"7E",X"01",X"FE",X"4C",X"DA",X"F4",X"0D",X"3A",X"15",X"90",X"A7",X"CA",X"F4",X"0D",
		X"3A",X"AD",X"92",X"A7",X"C2",X"F4",X"0D",X"EB",X"21",X"68",X"88",X"06",X"08",X"7E",X"FE",X"80",
		X"28",X"06",X"2C",X"2C",X"10",X"F7",X"18",X"6C",X"36",X"06",X"26",X"9B",X"36",X"01",X"E5",X"26",
		X"93",X"54",X"1D",X"1A",X"4F",X"77",X"1C",X"2C",X"1A",X"47",X"77",X"26",X"9B",X"54",X"1A",X"CB",
		X"0E",X"0F",X"CB",X"16",X"07",X"CB",X"18",X"3A",X"62",X"93",X"91",X"F5",X"30",X"02",X"ED",X"44",
		X"67",X"3A",X"15",X"92",X"A7",X"3E",X"95",X"28",X"02",X"3E",X"1C",X"90",X"30",X"02",X"ED",X"44",
		X"CD",X"A9",X"0E",X"44",X"4D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"09",X"CB",X"3C",
		X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"7C",X"A7",X"20",X"05",X"7D",X"FE",X"60",X"38",X"02",X"3E",
		X"60",X"47",X"F1",X"CB",X"18",X"E1",X"7D",X"C6",X"08",X"E6",X"0F",X"21",X"B0",X"92",X"85",X"6F",
		X"70",X"23",X"36",X"00",X"3A",X"E2",X"92",X"DD",X"77",X"0E",X"21",X"89",X"92",X"35",X"C8",X"11",
		X"14",X"00",X"DD",X"19",X"C3",X"E4",X"08",X"AF",X"DD",X"CB",X"13",X"86",X"DD",X"77",X"00",X"DD",
		X"77",X"02",X"26",X"88",X"DD",X"6E",X"10",X"36",X"02",X"26",X"8B",X"2C",X"7E",X"2D",X"3C",X"E6",
		X"07",X"FE",X"05",X"38",X"14",X"3A",X"2E",X"98",X"4F",X"E6",X"F8",X"C6",X"06",X"77",X"2C",X"79",
		X"E6",X"07",X"77",X"2D",X"3E",X"01",X"32",X"2D",X"98",X"DD",X"7E",X"06",X"DD",X"77",X"01",X"DD",
		X"7E",X"07",X"DD",X"77",X"03",X"C3",X"FE",X"0C",X"26",X"88",X"DD",X"6E",X"10",X"36",X"80",X"26",
		X"93",X"36",X"00",X"DD",X"36",X"13",X"00",X"C3",X"FA",X"0D",X"C5",X"D5",X"7B",X"95",X"06",X"00",
		X"30",X"04",X"CB",X"C0",X"ED",X"44",X"4F",X"7A",X"94",X"30",X"0A",X"57",X"78",X"EE",X"01",X"F6",
		X"02",X"47",X"7A",X"ED",X"44",X"B9",X"F5",X"17",X"A8",X"1F",X"3F",X"CB",X"10",X"F1",X"30",X"03",
		X"51",X"4F",X"7A",X"61",X"2E",X"00",X"CD",X"A9",X"0E",X"7C",X"A8",X"E6",X"01",X"28",X"03",X"7D",
		X"2F",X"6F",X"60",X"D1",X"C1",X"C9",X"D5",X"EB",X"21",X"00",X"00",X"CB",X"3F",X"30",X"01",X"19",
		X"CB",X"23",X"CB",X"12",X"A7",X"20",X"F4",X"D1",X"C9",X"C5",X"4F",X"AF",X"06",X"11",X"8F",X"38",
		X"0B",X"B9",X"38",X"01",X"91",X"3F",X"ED",X"6A",X"10",X"F4",X"C1",X"C9",X"91",X"37",X"C3",X"B6",
		X"0E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"06",X"68",X"E6",X"02",X"C0",
		X"21",X"FF",X"10",X"7E",X"2E",X"DF",X"4E",X"7E",X"A9",X"CB",X"67",X"20",X"01",X"C7",X"11",X"F7",
		X"89",X"21",X"F6",X"89",X"01",X"13",X"00",X"ED",X"B8",X"DD",X"21",X"D5",X"0F",X"1E",X"E0",X"01",
		X"04",X"05",X"DD",X"7E",X"00",X"DD",X"23",X"6F",X"26",X"10",X"7E",X"7B",X"81",X"5F",X"7E",X"12",
		X"10",X"F0",X"06",X"05",X"21",X"E4",X"89",X"7E",X"2C",X"B6",X"2C",X"2F",X"A6",X"2C",X"A6",X"2C",
		X"E6",X"0F",X"20",X"04",X"10",X"F1",X"18",X"40",X"05",X"28",X"4F",X"05",X"CB",X"20",X"CB",X"20",
		X"0F",X"38",X"03",X"04",X"18",X"FA",X"3A",X"E0",X"89",X"CB",X"3F",X"5F",X"CB",X"11",X"C6",X"E1",
		X"6F",X"26",X"89",X"7E",X"CB",X"41",X"28",X"04",X"07",X"07",X"07",X"07",X"E6",X"F0",X"B0",X"CB",
		X"41",X"28",X"04",X"07",X"07",X"07",X"07",X"77",X"3A",X"E0",X"89",X"A7",X"20",X"02",X"3E",X"02",
		X"3D",X"32",X"E0",X"89",X"7B",X"A7",X"28",X"09",X"2A",X"E2",X"89",X"7E",X"32",X"E1",X"89",X"18",
		X"42",X"2A",X"E2",X"89",X"3A",X"E1",X"89",X"77",X"18",X"39",X"4F",X"21",X"E0",X"89",X"CB",X"41",
		X"20",X"2D",X"7E",X"CB",X"3F",X"28",X"13",X"CB",X"59",X"20",X"0C",X"7E",X"FE",X"05",X"30",X"03",
		X"34",X"18",X"D5",X"36",X"05",X"18",X"D1",X"35",X"18",X"CE",X"2A",X"E2",X"89",X"CB",X"59",X"20",
		X"03",X"2B",X"18",X"01",X"23",X"22",X"E2",X"89",X"3E",X"01",X"32",X"E0",X"89",X"18",X"B9",X"36",
		X"05",X"18",X"B5",X"21",X"CA",X"83",X"11",X"E1",X"89",X"06",X"03",X"1A",X"1C",X"CD",X"C6",X"0F",
		X"10",X"F9",X"21",X"CA",X"87",X"3A",X"E0",X"89",X"06",X"06",X"A7",X"4F",X"28",X"02",X"0E",X"01",
		X"71",X"2C",X"3D",X"10",X"F5",X"C9",X"4F",X"E6",X"0F",X"77",X"2C",X"79",X"07",X"07",X"07",X"07",
		X"E6",X"0F",X"77",X"2C",X"C9",X"FD",X"FB",X"F7",X"EF",X"FE",X"23",X"00",X"1B",X"23",X"F0",X"40",
		X"23",X"00",X"09",X"23",X"05",X"11",X"23",X"00",X"10",X"23",X"10",X"40",X"23",X"04",X"30",X"FF",
		X"23",X"02",X"35",X"23",X"08",X"10",X"23",X"10",X"3C",X"23",X"00",X"FF",X"FF",X"AC",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
